LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY controller IS 
	PORT
	(
	CLR : IN STD_LOGIC;
	SWA : IN STD_LOGIC;
	SWB : IN STD_LOGIC;
	SWC : IN STD_LOGIC;
	IRH : IN STD_LOGIC_VECTOR (3 DOWNTO 0);
	C : IN STD_LOGIC;
	Z : IN STD_LOGIC;
	T3 : IN STD_LOGIC;
	W1 : IN STD_LOGIC;
	W2 : IN STD_LOGIC;
	W3 : IN STD_LOGIC;
	
	ABUS : OUT STD_LOGIC;
	ARINC : OUT STD_LOGIC;
	CIN : OUT STD_LOGIC;
	DRW : OUT STD_LOGIC;
	LAR : OUT STD_LOGIC;
	LDC : OUT STD_LOGIC;
	LDZ : OUT STD_LOGIC;
	LIR : OUT STD_LOGIC;
	LONG : OUT STD_LOGIC;
	LPC : OUT STD_LOGIC;
	M : OUT STD_LOGIC;
	MBUS : OUT STD_LOGIC;
	MEMW : OUT STD_LOGIC;
	PCADD : OUT STD_LOGIC;
	PCINC : OUT STD_LOGIC;
	S3 : OUT STD_LOGIC;
	S2 : OUT STD_LOGIC;
	S1 : OUT STD_LOGIC;
	S0 : OUT STD_LOGIC;
	SBUS : OUT STD_LOGIC;
	SEL3 : OUT STD_LOGIC;
	SEL2 : OUT STD_LOGIC;
	SEL1 : OUT STD_LOGIC;
	SEL0 : OUT STD_LOGIC;
	SELCTL : OUT STD_LOGIC;
	SHORT : OUT STD_LOGIC;
	STOP : OUT STD_LOGIC
	);
END controller;

ARCHITECTURE hardWireController of controller IS
	SIGNAL ST0, SST0, FLAG: STD_LOGIC;
BEGIN
	
	PROCESS(CLR, SWA, SWB, SWC, T3, IRH, W1, W2, W3, Z, C)
	VARIABLE WR : STD_LOGIC;
	VARIABLE RR : STD_LOGIC;
	VARIABLE WM : STD_LOGIC;
	VARIABLE RM : STD_LOGIC;
	VARIABLE EX : STD_LOGIC;
	VARIABLE SPC : STD_LOGIC;
	VARIABLE ADDI : STD_LOGIC;
	VARIABLE SUBI : STD_LOGIC;
	VARIABLE ANDI : STD_LOGIC;
	VARIABLE INCI : STD_LOGIC;
	VARIABLE LDI : STD_LOGIC;
	VARIABLE STI : STD_LOGIC;
	VARIABLE JCI : STD_LOGIC;
	VARIABLE JZI : STD_LOGIC;
	VARIABLE JMPI : STD_LOGIC;
	VARIABLE OUTI : STD_LOGIC;
	VARIABLE ORI : STD_LOGIC;
	VARIABLE DECI : STD_LOGIC;
	VARIABLE NOTI : STD_LOGIC;
	VARIABLE STPI : STD_LOGIC;
	VARIABLE NOPI : STD_LOGIC;
	BEGIN
	
	ABUS <= '0';
	ARINC <= '0';
	CIN <= '0';
	DRW <= '0';
	LAR <= '0';
	LDC <= '0';
	LDZ <= '0';
	LIR <= '0';
	LONG <= '0';
	LPC <= '0';
	M <= '0';
	MBUS <= '0';
	MEMW <= '0';
	PCADD <= '0';
	PCINC <= '0';
	S3 <= '0';
	S2 <= '0';
	S1 <= '0';
	S0 <= '0';
	SBUS <= '0';
	SEL3 <= '0';
	SEL2 <= '0';
	SEL1 <= '0';
	SEL0 <= '0';
	SELCTL <= '0';
	SHORT <= '0';
	STOP <= '0';
	
	ADDI := '0';
	SUBI := '0';
	ANDI := '0';
	INCI := '0';
	LDI := '0';
	STI := '0';
	JCI := '0';
	JZI := '0';
	JMPI := '0';
	OUTI := '0';
	ORI := '0';
	DECI := '0';
	NOTI := '0';
	STPI := '0';
	NOPI := '0';
	
	WR := SWC AND (NOT SWB) AND (NOT SWA);
	RR := (NOT SWC) AND SWB AND SWA;
	WM := (NOT SWC) AND (NOT SWB) AND SWA;
	RM := (NOT SWC) AND SWB AND (NOT SWA);
	
	IF (CLR = '0') THEN
		SST0 <= '0';
		ST0 <= '0';
		FLAG <= '0';
	ELSIF (T3'EVENT AND T3 = '0') THEN
		IF (SST0 = '1') THEN
			ST0 <= '1';
		ELSIF (WR = '1' AND FLAG = '1') THEN
			ST0 <= '0';
		END IF;
	END IF;
	
	IF (WR = '1' AND W2 = '1' AND ST0 = '1') THEN
		FLAG <= '1';
	ELSE 
		FLAG <= '0';
	END IF;
	
	EX := (NOT (SWC OR SWB OR SWA)) AND ST0;
	SPC := (NOT (SWC OR SWB OR SWA OR ST0));
	
	CASE IRH IS
		WHEN "0000" => NOPI := '1';
		WHEN "0001" => ADDI := '1';
		WHEN "0010" => SUBI := '1';
		WHEN "0011" => ANDI := '1';
		WHEN "0100" => INCI := '1';
		WHEN "0101" => LDI := '1';
		WHEN "0110" => STI := '1';
		WHEN "0111" => JCI := '1';
		WHEN "1000" => JZI := '1';
		WHEN "1001" => JMPI := '1';
		WHEN "1010" => OUTI := '1';
		WHEN "1011" => ORI := '1';
		WHEN "1100" => DECI := '1';
		WHEN "1101" => NOTI := '1';
		WHEN "1110" => STPI := '1';
		WHEN OTHERS => NOPI := '0';
	END CASE;
	
	ABUS <= (EX OR SPC) AND ((W2 AND (ADDI OR SUBI OR ANDI OR INCI OR LDI OR STI OR JMPI OR OUTI OR ORI OR DECI OR NOTI)) OR (W3 AND STI));
	ARINC <= ST0 AND W1 AND (RM OR WM);
	CIN <= (EX OR SPC) AND (W2 AND (ADDI OR DECI));
	DRW <= ((W1 OR W2) AND WR) OR ((EX OR SPC) AND ((W2 AND (ADDI OR SUBI OR ANDI OR INCI OR ORI OR DECI OR NOTI)) OR (W3 AND LDI)));
	LAR <= ((NOT ST0) AND W1 AND (RM OR WM)) OR ((EX OR SPC) AND (W2 AND (LDI OR STI)));
	LDC <= (EX OR SPC) AND (W2 AND (ADDI OR SUBI OR INCI OR DECI));
	LDZ <= (EX OR SPC) AND (W2 AND (ADDI OR SUBI OR ANDI OR INCI OR ORI OR DECI OR NOTI));
	LIR <= (EX) AND (NOT SPC) AND (W1 AND (ADDI OR SUBI OR ANDI OR INCI OR LDI OR STI OR JCI OR JZI OR JMPI OR OUTI OR ORI OR DECI OR NOTI OR STPI OR NOPI));
	LONG <= (EX OR SPC) AND (W2 AND (LDI OR STI));
	LPC <= ((NOT ST0) AND W1 AND SPC) OR ((EX OR SPC) AND (W2 AND JMPI));
	M <= (EX OR SPC) AND ((W2 AND (ANDI OR LDI OR STI OR JMPI OR ORI OR NOTI)) OR (W3 AND STI));
	MBUS <= (ST0 AND W1 AND RM) OR ((EX OR SPC) AND (W3 AND LDI));
	MEMW <= (ST0 AND W1 AND WM) OR ((EX OR SPC) AND (W3 AND STI));
	PCADD <= (EX OR SPC) AND ((C AND W2 AND JCI) OR (Z AND W2 AND JZI));
	PCINC <= (EX) AND (NOT SPC) AND (W1 AND (ADDI OR SUBI OR ANDI OR INCI OR LDI OR STI OR JCI OR JZI OR JMPI OR OUTI OR ORI OR DECI OR NOTI OR STPI OR NOPI));
	S3 <= (EX OR SPC) AND ((W2 AND (ADDI OR ANDI OR LDI OR STI OR JMPI OR OUTI OR ORI OR DECI)) OR (W3 AND STI));
	S2 <= (EX OR SPC) AND (W2 AND (SUBI OR (W2 AND STI) OR JMPI OR ORI OR DECI));
	S1 <= (EX OR SPC) AND ((W2 AND (SUBI OR ANDI OR LDI OR STI OR JMPI OR OUTI OR ORI OR DECI)) OR (W3 AND STI));
	S0 <= (EX OR SPC) AND (W2 AND (ADDI OR ANDI OR (W2 AND STI) OR JMPI OR DECI));
	SBUS <= ((NOT ST0) AND W1 AND (RM OR SPC)) OR (W1 AND (WM OR WR)) OR (W2 AND WR);
	SEL3 <= (ST0 AND WR AND (W1 OR W2)) OR (W2 AND RR);
	SEL2 <= W2 AND WR;
	SEL1 <= (((NOT ST0 AND W1) OR (ST0 AND W2)) AND WR) OR (W2 AND RR);
	SEL0 <= (W1 AND (RR OR WR)) OR (W2 AND RR);
	SELCTL <= ((W1 OR W2) AND (RR OR WR)) OR (W1 AND (RM OR WM)) OR ((NOT ST0) AND W1 AND SPC);
	SHORT <= (W1 AND (RM OR WM)) OR ((NOT ST0) AND W1 AND SPC);
	STOP <= ((W1 OR W2) AND (WR OR RR)) OR (W1 AND (RM OR WM)) OR ((NOT ST0) AND W1 AND SPC) OR ((EX OR SPC) AND W2 AND STPI);
	SST0 <= (W2 AND WR AND (NOT ST0)) OR (W1 AND (RM OR WM) AND (NOT ST0)) OR ((NOT ST0) AND W1 AND SPC);	

	END PROCESS;
END ARCHITECTURE;
